interface intf(input logic clk, reset);
    logic [7:0] in_a, in_b;
    logic [8:0] out;
  endinterface
